** Profile: "SCHEMATIC1-potectie_temperatura"  [ c:\users\bianca\desktop\p1_2023_431e_naftanaila_bianca_elena_sers_n16_orcad\schematics\stabilizator de tensiune cu ers\stabilizator_de_tensiune_ers-pspicefiles\schematic1\potectie_temperatura.sim ] 

** Creating circuit file "potectie_temperatura.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "c:/users/bianca/desktop/modele_leduri/smls14bet.lib" 
.LIB "c:/users/bianca/desktop/modele_a1_lib/bc807-25.lib" 
.LIB "c:/users/bianca/desktop/modele_a1_lib/bc817-25.lib" 
.LIB "c:/users/bianca/desktop/modele_a1_lib/bc846b.lib" 
.LIB "c:/users/bianca/desktop/modele_a1_lib/bzx84c2v7.lib" 
.LIB "c:/users/bianca/desktop/modele_a1_lib/bzx84c5v1.lib" 
.LIB "c:/users/bianca/desktop/modele_a1_lib/mjd31cg.lib" 
* From [PSPICE NETLIST] section of C:\Users\Bianca\AppData\Local\Temp\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC LIN TEMP -20 120 1 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
